----------------------------------------------------------------------
-- Fichero: MicroSuma.vhd
-- Descripci�n:
-- Fecha �ltima modificaci�n: 2016-02-24

-- Autores: Jos� Ignacio G�mez (2016), �scar G�mez (2016) 
-- Asignatura: E.C. 1� grado
-- Grupo de Pr�cticas: 2101
-- Grupo de Teor�a:210
-- Pr�ctica: 2
-- Ejercicio: 2
----------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.std_LOGIC_arith.ALL;
use IEEE.std_logic_unsigned.ALL;

